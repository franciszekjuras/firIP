
`timescale 1 ns / 1 ps

	module firMainAXI #
	(
		// Users to add parameters here
		parameter FIR_DATA_WIDTH = 14,
		parameter FIR_COEF_WIDTH = 18,
		parameter FIR_COEF_MAG = 0,
		parameter FIR_DSP_NR = 4, 
		parameter FIR_TM = 2,

		// User parmaters end

		parameter integer C_S_AXI_DATA_WIDTH	= 32,
		parameter integer C_S_AXI_ADDR_WIDTH	= 16
	)
	(
		// Users to add ports here
		input wire fir_clk,
		input wire signed [FIR_DATA_WIDTH-1 : 0] fir_in,
		output reg signed [FIR_DATA_WIDTH-1 : 0] fir_out,
		output wire [7:0] leds_out,
		// User ports ends
		
		input wire  S_AXI_ACLK,
		input wire  S_AXI_ARESETN,
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_AWADDR,
		input wire [2 : 0] S_AXI_AWPROT,
		input wire  S_AXI_AWVALID,
		output wire  S_AXI_AWREADY,
		input wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_WDATA,
		input wire [(C_S_AXI_DATA_WIDTH/8)-1 : 0] S_AXI_WSTRB,
		input wire  S_AXI_WVALID,
		output wire  S_AXI_WREADY,
		output wire [1 : 0] S_AXI_BRESP,
		output wire  S_AXI_BVALID,
		input wire  S_AXI_BREADY,
		input wire [C_S_AXI_ADDR_WIDTH-1 : 0] S_AXI_ARADDR,
		input wire [2 : 0] S_AXI_ARPROT,
		input wire  S_AXI_ARVALID,
		output wire  S_AXI_ARREADY,
		output wire [C_S_AXI_DATA_WIDTH-1 : 0] S_AXI_RDATA,
		output wire [1 : 0] S_AXI_RRESP,
		output wire  S_AXI_RVALID,
		input wire  S_AXI_RREADY
	);
	
	// local parameter for addressing 32 bit / 64 bit C_S_AXI_DATA_WIDTH
	// ADDR_LSB is used for addressing 32/64 bit registers/memories
	// ADDR_LSB = 2 for 32 bits addressing
	// ADDR_LSB = 3 for 64 bits addressing

	localparam FIR_COEFS_NR = FIR_TM * FIR_DSP_NR;

	localparam ADDR_LSB = (C_S_AXI_DATA_WIDTH/32) + 1;
	// Addresses' bases in 32/64 bit addressing
	localparam FIR_OFFSET_COEFS = 8;
	localparam FIR_OFFSET_DEBUG = 128;
	//reverse order xD
	localparam PROG_NAME = "_RIF";
	localparam PROG_VER = "2MT";

	//Switches:
	localparam SWITCH_CON_EST = 0;
	localparam SWITCH_FIR_EN = 1;
	localparam SWITCH_FIR_UPDATE = 2;
	localparam SWITCH_FIR_SNAP = 5;
	localparam SWITCH_FIR_DEBUG_1 = 6;
	localparam SWITCH_FIR_DEBUG_2 = 7;
	//Debug switches:

	integer idx;

	// AXI4LITE signals
	reg [C_S_AXI_ADDR_WIDTH - ADDR_LSB -1 : 0] 	axi_awaddr;
	reg  	axi_awready;
	reg  	axi_wready;
	reg [1 : 0] 	axi_bresp;
	reg  	axi_bvalid;
	reg [C_S_AXI_ADDR_WIDTH - ADDR_LSB -1 : 0] 	axi_araddr;
	reg  	axi_arready;
	reg [C_S_AXI_DATA_WIDTH-1 : 0] 	axi_rdata;
	reg [1 : 0] 	axi_rresp;
	reg  	axi_rvalid;
	wire	 reg_rden;
	wire	 reg_wren;
	reg [C_S_AXI_DATA_WIDTH-1:0]	 reg_data_out;
	reg	 aw_en;

	// I/O Connections assignments
	assign S_AXI_AWREADY	= axi_awready;
	assign S_AXI_WREADY	= axi_wready;
	assign S_AXI_BRESP	= axi_bresp;
	assign S_AXI_BVALID	= axi_bvalid;
	assign S_AXI_ARREADY	= axi_arready;
	assign S_AXI_RDATA	= axi_rdata;
	assign S_AXI_RRESP	= axi_rresp;
	assign S_AXI_RVALID	= axi_rvalid;

	// Registers connected to AXI
	//read-only
/*0*/    reg [C_S_AXI_DATA_WIDTH-1 : 0] info_1;
/*1*/    reg [C_S_AXI_DATA_WIDTH-1 : 0] info_2; //TODO: add extra info,
/*2*/    reg [C_S_AXI_DATA_WIDTH-1 : 0] coefs_max_nr;
/*3*/    //reg [C_S_AXI_DATA_WIDTH-1 : 0] unused;
	//write|read
/*4*/    reg [C_S_AXI_DATA_WIDTH-1 : 0] switches;
/*5*/    reg [C_S_AXI_DATA_WIDTH-1 : 0] coefs_crr_nr;
/*6*/    //reg [C_S_AXI_DATA_WIDTH-1 : 0] unused;
/*7*/    //reg [C_S_AXI_DATA_WIDTH-1 : 0] unused;

	reg signed [FIR_COEF_WIDTH-1 : 0] coefs [FIR_COEFS_NR];

	/*Dozen of boring AXI4-lite procedures*/
	always @( posedge S_AXI_ACLK ) begin
	if ( S_AXI_ARESETN == 1'b0 ) begin
		axi_awready <= 1'b0;
		aw_en <= 1'b1;
		end else begin    
		if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en) begin
			axi_awready <= 1'b1;
			aw_en <= 1'b0;
			end else if (S_AXI_BREADY && axi_bvalid) begin
				aw_en <= 1'b1;
				axi_awready <= 1'b0;
			end else begin
				axi_awready <= 1'b0;
			end
		end 
	end       

	always @( posedge S_AXI_ACLK )begin
		if ( S_AXI_ARESETN == 1'b0 )
			axi_awaddr <= 0;
		else begin    
			if (~axi_awready && S_AXI_AWVALID && S_AXI_WVALID && aw_en)
				axi_awaddr <= S_AXI_AWADDR[C_S_AXI_ADDR_WIDTH-1 : ADDR_LSB];
		end 
	end       

	always @( posedge S_AXI_ACLK )begin
		if ( S_AXI_ARESETN == 1'b0 )
			axi_wready <= 1'b0;
		else begin    
			if (~axi_wready && S_AXI_WVALID && S_AXI_AWVALID && aw_en) 
				axi_wready <= 1'b1;
			else
				axi_wready <= 1'b0;
		end 
	end       

	assign reg_wren = axi_wready && S_AXI_WVALID && axi_awready && S_AXI_AWVALID;

	//-----------------------------------------------------//
	//--------------------WRITE MAPPING--------------------//
	//-----------------------------------------------------//

	always @( posedge S_AXI_ACLK ) begin: write_data
		if (reg_wren & S_AXI_ARESETN) begin
			for(idx = 0; idx < FIR_COEFS_NR; idx = idx + 1) begin
				if(idx + FIR_OFFSET_COEFS == axi_awaddr)
					coefs[idx] <= {S_AXI_WDATA[C_S_AXI_DATA_WIDTH-1],S_AXI_WDATA[FIR_COEF_WIDTH-2 : 0]};
			end

			case(axi_awaddr)
				4: switches <= S_AXI_WDATA;
				5: coefs_crr_nr <= S_AXI_WDATA;
				//6: unused <= S_AXI_WDATA;
				//7: unused <= S_AXI_WDATA;
			endcase
		end
	end    

	always @( posedge S_AXI_ACLK ) begin
		if ( S_AXI_ARESETN == 1'b0 ) begin
			axi_bvalid  <= 0;
			axi_bresp   <= 2'b0;
		end else begin    
			if (axi_awready && S_AXI_AWVALID && ~axi_bvalid && axi_wready && S_AXI_WVALID) begin
				axi_bvalid <= 1'b1;
				axi_bresp  <= 2'b0; // 'OKAY' response 
			end else begin
				if (S_AXI_BREADY && axi_bvalid)
					axi_bvalid <= 1'b0; 
			end
		end
	end   

	always @( posedge S_AXI_ACLK ) begin
		if ( S_AXI_ARESETN == 1'b0 ) begin
			axi_arready <= 1'b0;
			axi_araddr  <= 32'b0;
		end else begin    
			if (~axi_arready && S_AXI_ARVALID) begin
				axi_arready <= 1'b1;
				axi_araddr  <= S_AXI_ARADDR[C_S_AXI_ADDR_WIDTH-1 : ADDR_LSB];
			end else begin
				axi_arready <= 1'b0;
			end
		end 
	end

	always @( posedge S_AXI_ACLK ) begin
		if ( S_AXI_ARESETN == 1'b0 ) begin
			axi_rvalid <= 0;
			axi_rresp  <= 0;
		end else begin    
			if (axi_arready && S_AXI_ARVALID && ~axi_rvalid) begin
				axi_rvalid <= 1'b1;
				axi_rresp  <= 2'b0; // 'OKAY' response
			end else if (axi_rvalid && S_AXI_RREADY) begin
			  axi_rvalid <= 1'b0;
			end                
		end
	end 

	//-----------------------------------------------------//
	//---------------------READ MAPPING--------------------//
	//-----------------------------------------------------//

	assign reg_rden = axi_arready & S_AXI_ARVALID & ~axi_rvalid;
	always @(*)
	begin
		// Address decoding for reading registers
		case ( axi_araddr )
		0 : reg_data_out = info_1;
		1 : reg_data_out = info_2;
		2 : reg_data_out = coefs_max_nr;
		// 3 : reg_data_out = unused;
		4 : reg_data_out = switches;
		5 : reg_data_out = coefs_crr_nr;
		// 6 : reg_data_out = unused;
		// 7 : reg_data_out = unused;
		default : reg_data_out = 0;
		endcase
		/*IF COEFS STATUS IS NECESSARY*/
		for(idx = 0; idx < (DEBUG_LENGTH*DEBUG_DEPTH); idx = idx + 1) begin
			if(idx + FIR_OFFSET_DEBUG == axi_araddr) begin
				reg_data_out = debug_block[idx]; //WARN:sign bit might not be shifted properly
			end
		end	   
	end

	always @( posedge S_AXI_ACLK ) begin
		if ( S_AXI_ARESETN == 1'b0 ) begin
			axi_rdata  <= 0;
		end else begin 
			if (reg_rden)
				axi_rdata <= reg_data_out;
		end
	end    

	//-----------------------------------------------------//
	//------------------------LOGIC------------------------//
	//-----------------------------------------------------//

	//LEDS
	assign leds_out[7:0] = switches[7:0];

	//COUNTER
	localparam COUNT_WIDTH = $clog2(FIR_TM);
	wire [COUNT_WIDTH-1:0] count;

	counter #(
	.COUNT_WIDTH(COUNT_WIDTH),
	.MODULO(FIR_TM)) 
	inst_counter (
	.clk(fir_clk),
	.count(count));

	//counter connections wiring
	wire [COUNT_WIDTH-1:0] dsp_con_count [FIR_DSP_NR + 1];
	assign dsp_con_count[0] = count;
	// localparam DSP_MULT_LAT_DIFF = 1; // latency difference between coef and sample input
	// shiftby #(.BY(DSP_MULT_LAT_DIFF), .WIDTH(COUNT_WIDTH))
	// shift_coef_count 
	// (.in(count), .out(dsp_con_count[0]), .clk(fir_clk));



	localparam SUM_WIDTH = FIR_DATA_WIDTH + FIR_COEF_MAG; /*at the end, sum is shortened by COEFMAG to XW length,
	so there is little reason to add more registers*/

	wire signed [SUM_WIDTH-1:0] dsp_con_sum [FIR_DSP_NR:0]; //+1 because of beg and end, ex: ---DSP---DSP---DSP--- || note: 3 DSPs and 4 wires
	wire signed [FIR_DATA_WIDTH-1:0] dsp_con_x [FIR_DSP_NR:0]; //same as above
	
	wire signed [SUM_WIDTH-1:0] sum_loop_end;
	wire signed [FIR_DATA_WIDTH-1:0] data_loop_end;
	localparam LOOP_FEEDBACK_SYNC = FIR_TM + 1 - (FIR_DSP_NR%FIR_TM);

	shiftby #(.BY(LOOP_FEEDBACK_SYNC), .WIDTH(SUM_WIDTH))
	shift_data_loop
	(.in(dsp_con_x[FIR_DSP_NR]), .out(data_loop_end), .clk(fir_clk));

	shiftby #(.BY(LOOP_FEEDBACK_SYNC), .WIDTH(FIR_DATA_WIDTH))
	shift_sum_loop
	(.in(dsp_con_sum[FIR_DSP_NR]), .out(sum_loop_end), .clk(fir_clk));


	loop_multplx #(
	.COUNT_WIDTH(COUNT_WIDTH),
	.DATA_WIDTH(FIR_DATA_WIDTH)	
	) 
	inst_in_multplx (
	.count(count),
	.in(fir_in),
	.loop(data_loop_end),
	.out(dsp_con_x[0])
	);


	localparam DSP_PIPELINE_DIFF = 1; // difference in registers from in multiplexers to first summation in dsp block (so fresh sample would contribute to fresh 0 sum)
	wire [COUNT_WIDTH-1:0] sum_count;
	shiftby #(.BY(DSP_PIPELINE_DIFF), .WIDTH(COUNT_WIDTH))
	shift_sum_count 
	(.in(count), .out(sum_count), .clk(fir_clk));

	loop_multplx #(
	.COUNT_WIDTH(COUNT_WIDTH),
	.DATA_WIDTH(FIR_DATA_WIDTH)	
	) 
	inst_sum_multplx (
	.count(sum_count),
	.in(0),
	.loop(sum_loop_end),
	.out(dsp_con_sum[0])
	);

	// always @(posedge fir_clk) begin
	// 	if(switches[SWITCH_FIR_EN] == 1'b1) begin
	// 		fir_out[FIR_DATA_WIDTH-1:0] <= dsp_con_sum[FIR_DSP_NR][SUM_WIDTH-1: SUM_WIDTH - FIR_DATA_WIDTH]; 
	// 		//output shift by coefficients' magnitude
	// 		//same as [FIR_COEF_MAG + FIR_DATA_WIDTH - 1 : FIR_COEF_MAG] 
	// 	end else begin
	// 		fir_out <= fir_in;
	// 	end
	// end
	// Generating fir taps (DSP blocks + shifting registers + coefficients' multiplexers)
		//coef_mult wiring

	reg signed [FIR_COEF_WIDTH-1 : 0] coefs_pack [FIR_DSP_NR][FIR_TM];
	genvar i_cp, j_cp;
	for(i_cp = 0; i_cp < FIR_DSP_NR; i_cp = i_cp + 1) begin
		for(j_cp = 0; j_cp < FIR_TM; j_cp = j_cp + 1) begin
			assign coefs_pack[i_cp][j_cp] = coefs[FIR_DSP_NR * j_cp + i_cp];
		end
	end


	wire signed [FIR_COEF_WIDTH-1 : 0] coef_crr [FIR_DSP_NR];

	wire signed [FIR_COEF_WIDTH-1 : 0] coef_crr_debug1 [FIR_DSP_NR];
	reg signed [FIR_COEF_WIDTH-1 : 0] coef_crr_debug2 [FIR_DSP_NR];

	generate
		for(genvar k = 0; k < FIR_DSP_NR; k = k + 1) begin
			firtap #(
			.XW(FIR_DATA_WIDTH),
			.COEFW(FIR_COEF_WIDTH),
			.OUTW(SUM_WIDTH),
			.SAMPLE_SHIFT(1),
			.SUM_SHIFT(1+FIR_TM)
			) inst_tap(
			.clk(fir_clk),
			.inX(dsp_con_x[k]),
			.outX(dsp_con_x[k+1]),
			.inCoef(coef_crr[k]),
			.inSum(dsp_con_sum[k]),
			.outSum(dsp_con_sum[k+1])
			);
		end
	endgenerate

	generate
		for(genvar l = 0; l < FIR_DSP_NR; l = l+1) begin
			coef_multplx #(
			.COEFW(FIR_COEF_WIDTH),
			.TM(FIR_TM),
			.CW(COUNT_WIDTH)
			) inst_coef_multplx(
			.clk(fir_clk),
			.counter_in(dsp_con_count[l]),
			.counter_out(dsp_con_count[l+1]),
			.coef_pack(coefs_pack[l]),
			.coef_out(coef_crr[l])
			);
		end
	endgenerate
	// generate		
	// 	for(genvar k = 0; k < FIR_DSP_NR; k = k + 1) begin
	// 		coef_multplx #(
	// 		.COEFW(FIR_COEF_WIDTH),
	// 		.TM(FIR_TM),
	// 		.CW(COUNT_WIDTH)
	// 		) inst_coef_multplx(
	// 		.clk(fir_clk),
	// 		.counter_in(dsp_con_count[k]),
	// 		.counter_out(dsp_con_count[k+1]),
	// 		.coef_pack(coefs_pack[k]),
	// 		.coef_out(coef_crr[k])
	// 		);
	// 	end
	// endgenerate

	// generate
	// 	for(genvar l = 0; k < FIR_DSP_NR; k = k + 1) begin
	// 		assign coef_crr_debug1[k] = coefs_pack[k][dsp_con_count[k]];
	// 	end
	// endgenerate
	// reg[31:0] cidx;
	// generate
	// 	for(genvar m = 0; k < FIR_DSP_NR; k = k + 1) begin
	// 		always_comb begin
	// 			for(cidx = 0; cidx < FIR_TM; cidx = cidx + 1)
	// 			begin
	// 				if(dsp_con_count[k] == cidx)
	// 					coef_crr_debug2[k] = 1024;
	// 			end
	// 		end
	// 	end
	// endgenerate




	//out
	reg [FIR_DATA_WIDTH-1:0] fir_in_debug_1;
	reg [FIR_DATA_WIDTH-1:0] fir_in_debug_2;
	reg [FIR_DATA_WIDTH-1:0]fir_in_debug_3;
	reg signed [FIR_DATA_WIDTH-1:0]sum_loop_out;
	reg [SUM_WIDTH-1:0]sum_loop_out_debug;
	always @(posedge fir_clk) begin
		if(sum_count == 0)
			sum_loop_out[FIR_DATA_WIDTH-1:0] <= sum_loop_end[SUM_WIDTH-1: SUM_WIDTH - FIR_DATA_WIDTH];
	end
	always @(posedge fir_clk) begin
		if(sum_count == 0)
			sum_loop_out_debug <= sum_loop_end;
	end
	always @(posedge fir_clk) begin
		fir_in_debug_3 <= fir_in;
	end
	always @(posedge fir_clk) begin
		if(count == 0) begin
			fir_in_debug_1 <= fir_in;
			fir_in_debug_2 <= fir_in;			
		end else begin
			fir_in_debug_2 <= 0;
		end
	end

	always @(*)
	begin
		case ({switches[SWITCH_FIR_EN],switches[SWITCH_FIR_DEBUG_1],switches[SWITCH_FIR_DEBUG_2]})
			3'b000	:	fir_out = fir_in;
			3'b100	:	fir_out = sum_loop_out;
			default	:	fir_out = 4096;
		endcase
	end

	assign debug1_in = dsp_con_sum[0];
	assign debug2_in = dsp_con_x[0];
	assign debug3_in = coef_crr[0];
	assign debug4_in = dsp_con_sum[1];
	assign debug5_in = dsp_con_x[1];
	assign debug6_in = coef_crr[1];
	assign debug7_in = dsp_con_sum[2];
	assign debug8_in = dsp_con_x[2];
	assign debug9_in = coef_crr[2];
	assign debug10_in = dsp_con_sum[3];


	/////////////////////

	always @(*) begin
		coefs_max_nr = FIR_COEFS_NR;
		info_1 = PROG_NAME;
		info_2 = PROG_VER; 
	end
	// User logic ends

	localparam DEBUG_LENGTH = 64;
	localparam DEBUG_DEPTH = 10;

	///////////////////////
	wire [C_S_AXI_DATA_WIDTH-1:0] debug1_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug1 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug1[0] <= debug1_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug1[k] <= debug1[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug2_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug2 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug2[0] <= debug2_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug2[k] <= debug2[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug3_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug3 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug3[0] <= debug3_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug3[k] <= debug3[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug4_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug4 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug4[0] <= debug4_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug4[k] <= debug4[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug5_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug5 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug5[0] <= debug5_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug5[k] <= debug5[k-1];
	        end
	    end
	end


	wire [C_S_AXI_DATA_WIDTH-1:0] debug6_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug6 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug6[0] <= debug6_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug6[k] <= debug6[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug7_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug7 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug7[0] <= debug7_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug7[k] <= debug7[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug8_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug8 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug8[0] <= debug8_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug8[k] <= debug8[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug9_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug9 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug9[0] <= debug9_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug9[k] <= debug9[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug10_in;
	reg [C_S_AXI_DATA_WIDTH-1:0] debug10 [DEBUG_LENGTH];
	integer k;
	always @(posedge fir_clk)
	begin
		if(switches[SWITCH_FIR_SNAP])
		begin
			debug10[0] <= debug10_in;
			for(k = 1; k < DEBUG_LENGTH; k = k + 1) begin
	            debug10[k] <= debug10[k-1];
	        end
	    end
	end

	wire [C_S_AXI_DATA_WIDTH-1:0] debug_block [DEBUG_LENGTH*DEBUG_DEPTH];
	genvar ideb;
	generate
		for(ideb = 0; ideb < DEBUG_LENGTH; ideb = ideb + 1) begin
			assign debug_block[ideb+(DEBUG_LENGTH*0)] = debug1[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*1)] = debug2[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*2)] = debug3[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*3)] = debug4[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*4)] = debug5[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*5)] = debug6[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*6)] = debug7[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*7)] = debug8[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*8)] = debug9[ideb];
			assign debug_block[ideb+(DEBUG_LENGTH*9)] = debug10[ideb];
		end
	endgenerate

	endmodule